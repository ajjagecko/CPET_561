
module nios_system (
	clk_clk,
	leds_export,
	pushbutton1_export);	

	input		clk_clk;
	output	[7:0]	leds_export;
	input		pushbutton1_export;
endmodule
